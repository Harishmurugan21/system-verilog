class transaction;
  rand logic[2:0] a;
  rand bit b;
  
endclass
  
 
