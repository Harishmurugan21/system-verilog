# transaction object get fro  driver a=000,b=0
# transaction object get fro  driver a=001,b=0
# transaction object get fro  driver a=100,b=1
# transaction object get fro  driver a=100,b=0
# transaction object get fro  driver a=111,b=1
