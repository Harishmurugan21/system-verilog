Compiler version U-2023.03-SP2_Full64; Runtime version U-2023.03-SP2_Full64;  Dec 16 13:04 2025
generator class signal
a=1,b=1,c=1,sum=0,carry=0
generator class signal
a=1,b=0,c=1,sum=0,carry=0
generator class signal
a=1,b=1,c=1,sum=0,carry=0
generator class signal
a=0,b=0,c=1,sum=0,carry=0
generator class signal
a=0,b=1,c=1,sum=0,carry=0
generator class signal
a=1,b=0,c=0,sum=0,carry=0
generator class signal
a=0,b=1,c=1,sum=0,carry=0
generator class signal
a=0,b=1,c=1,sum=0,carry=0
generator class signal
a=1,b=1,c=1,sum=0,carry=0
generator class signal
a=1,b=1,c=1,sum=0,carry=0
generator class signal
a=0,b=0,c=1,sum=0,carry=0
generator class signal
a=0,b=0,c=0,sum=0,carry=0
generator class signal
a=1,b=1,c=0,sum=0,carry=0
generator class signal
a=1,b=1,c=1,sum=0,carry=0
generator class signal
a=0,b=1,c=1,sum=0,carry=0
driver signal
a=1,b=1,c=1,sum=0,carry=0
monitor class signals
a=1,b=1,c=1,sum=1,carry=1
signals received on score board
a=1,b=1,c=1,sum=1,carry=1
--------pass-------
driver signal
a=1,b=0,c=1,sum=0,carry=0
monitor class signals
a=1,b=0,c=1,sum=0,carry=1
signals received on score board
a=1,b=0,c=1,sum=0,carry=1
--------pass-------
driver signal
a=1,b=1,c=1,sum=0,carry=0
monitor class signals
a=1,b=1,c=1,sum=1,carry=1
signals received on score board
a=1,b=1,c=1,sum=1,carry=1
--------pass-------
driver signal
a=0,b=0,c=1,sum=0,carry=0
monitor class signals
a=0,b=0,c=1,sum=1,carry=0
signals received on score board
a=0,b=0,c=1,sum=1,carry=0
--------pass-------
driver signal
a=0,b=1,c=1,sum=0,carry=0
monitor class signals
a=0,b=1,c=1,sum=0,carry=1
signals received on score board
a=0,b=1,c=1,sum=0,carry=1
--------pass-------
driver signal
a=1,b=0,c=0,sum=0,carry=0
monitor class signals
a=1,b=0,c=0,sum=1,carry=0
signals received on score board
a=1,b=0,c=0,sum=1,carry=0
--------pass-------
driver signal
a=0,b=1,c=1,sum=0,carry=0
monitor class signals
a=0,b=1,c=1,sum=0,carry=1
signals received on score board
a=0,b=1,c=1,sum=0,carry=1
--------pass-------
driver signal
a=0,b=1,c=1,sum=0,carry=0
monitor class signals
a=0,b=1,c=1,sum=0,carry=1
signals received on score board
a=0,b=1,c=1,sum=0,carry=1
--------pass-------
driver signal
a=1,b=1,c=1,sum=0,carry=0
monitor class signals
a=1,b=1,c=1,sum=1,carry=1
signals received on score board
a=1,b=1,c=1,sum=1,carry=1
--------pass-------
driver signal
a=1,b=1,c=1,sum=0,carry=0
monitor class signals
a=1,b=1,c=1,sum=1,carry=1
signals received on score board
a=1,b=1,c=1,sum=1,carry=1
--------pass-------
driver signal
a=0,b=0,c=1,sum=0,carry=0
monitor class signals
a=0,b=0,c=1,sum=1,carry=0
signals received on score board
a=0,b=0,c=1,sum=1,carry=0
--------pass-------
driver signal
a=0,b=0,c=0,sum=0,carry=0
monitor class signals
a=0,b=0,c=0,sum=0,carry=0
signals received on score board
a=0,b=0,c=0,sum=0,carry=0
--------pass-------
driver signal
a=1,b=1,c=0,sum=0,carry=0
monitor class signals
a=1,b=1,c=0,sum=0,carry=1
signals received on score board
a=1,b=1,c=0,sum=0,carry=1
--------pass-------
driver signal
a=1,b=1,c=1,sum=0,carry=0
monitor class signals
a=1,b=1,c=1,sum=1,carry=1
signals received on score board
a=1,b=1,c=1,sum=1,carry=1
--------pass-------
driver signal
a=0,b=1,c=1,sum=0,carry=0
monitor class signals
a=0,b=1,c=1,sum=0,carry=1
signals received on score board
a=0,b=1,c=1,sum=0,carry=1
--------pass-------
$finish at simulation time 
